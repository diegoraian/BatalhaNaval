module geracaoAleatoria (
    input clock,
    input reset,
    output [12:0] rnd
    );
	
	reg[3:0] x =3'd00;
	
 
endmodule