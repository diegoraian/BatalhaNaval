/*******************************************************************************

-- File Type:    Verilog HDL 
-- Tool Version: VHDL2verilog 20.20
-- Input file was: ..\..\..\..\OneDrive\1 - UFBA 5 semestre mexer aquiii\ENGG52 - Lab Integrado 1\PARA A ATIVIDADE 2\ARQUIVOS CONVERTIDOS EMBARCADOS ASCII\lista_caracteres_asteriscos\lista_caracteres_asteriscos_ece320web.vhd
-- Command line was: D:\SynaptiCAD\bin\win32\vhdl2verilog.exe ..\..\..\..\OneDrive\1 - UFBA 5 semestre mexer aquiii\ENGG52 - Lab Integrado 1\PARA A ATIVIDADE 2\ARQUIVOS CONVERTIDOS EMBARCADOS ASCII\lista_caracteres_asteriscos\lista_caracteres_asteriscos_ece320web.vhd -ncc
-- Date Created: Sun Aug 06 16:28:26 2017

*******************************************************************************/

`define false 1'b 0
`define FALSE 1'b 0
`define true 1'b 1
`define TRUE 1'b 1

`timescale 1 ns / 1 ns // timescale for following modules


//  Listing 13.1
//  ROM with synchonous read (inferring Block RAM)
//  character ROM
//    - 8-by-16 (8-by-2^4) font
//    - 128 (2^7) characters
//    - ROM size: 512-by-8 (2^11-by-8) bits
//                16K bits: 1 BRAM

module font_rom (
   clk,
   addr,
   data);
 

input   clk; 
input   [10:0] addr; 
output   [7:0] data; 

wire    [7:0] data; 
parameter ADDR_WIDTH = 11; 
parameter DATA_WIDTH = 8; 
reg     [ADDR_WIDTH - 1:0] addr_reg; 

//  ROM definition
parameter [DATA_WIDTH - 1:0] ROM = {8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 01111110, 8'b 10000001, 8'b 10100101, 8'b 10000001, 8'b 10000001, 8'b 10111101, 8'b 10011001, 8'b 10000001, 8'b 10000001, 8'b 01111110, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 01111110, 8'b 11111111, 8'b 11011011, 8'b 11111111, 8'b 11111111, 8'b 11000011, 8'b 11100111, 8'b 11111111, 8'b 11111111, 8'b 01111110, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 01101100, 8'b 11111110, 8'b 11111110, 8'b 11111110, 8'b 11111110, 8'b 01111100, 8'b 00111000, 8'b 00010000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00010000, 8'b 00111000, 8'b 01111100, 8'b 11111110, 8'b 01111100, 8'b 00111000, 8'b 00010000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00011000, 8'b 00111100, 8'b 00111100, 8'b 11100111, 8'b 11100111, 8'b 11100111, 8'b 00011000, 8'b 00011000, 8'b 00111100, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00011000, 8'b 00111100, 8'b 01111110, 8'b 11111111, 8'b 11111111, 8'b 01111110, 8'b 00011000, 8'b 00011000, 8'b 00111100, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00011000, 8'b 00111100, 8'b 00111100, 8'b 00011000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 11111111, 8'b 11111111, 8'b 11111111, 8'b 11111111, 8'b 11111111, 8'b 11111111, 8'b 11100111, 8'b 11000011, 8'b 11000011, 8'b 11100111, 8'b 11111111, 8'b 11111111, 8'b 11111111, 8'b 11111111, 8'b 11111111, 8'b 11111111, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00111100, 8'b 01100110, 8'b 01000010, 8'b 01000010, 8'b 01100110, 8'b 00111100, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 11111111, 8'b 11111111, 8'b 11111111, 8'b 11111111, 8'b 11111111, 8'b 11000011, 8'b 10011001, 8'b 10111101, 8'b 10111101, 8'b 10011001, 8'b 11000011, 8'b 11111111, 8'b 11111111, 8'b 11111111, 8'b 11111111, 8'b 11111111, 8'b 00000000, 8'b 00000000, 8'b 00011110, 8'b 00001110, 8'b 00011010, 8'b 00110010, 8'b 01111000, 8'b 11001100, 8'b 11001100, 8'b 11001100, 8'b 11001100, 8'b 01111000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00111100, 8'b 01100110, 8'b 01100110, 8'b 01100110, 8'b 01100110, 8'b 00111100, 8'b 00011000, 8'b 01111110, 8'b 00011000, 8'b 00011000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00111111, 8'b 00110011, 8'b 00111111, 8'b 00110000, 8'b 00110000, 8'b 00110000, 8'b 00110000, 8'b 01110000, 8'b 11110000, 8'b 11100000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 01111111, 8'b 01100011, 8'b 01111111, 8'b 01100011, 8'b 01100011, 8'b 01100011, 8'b 01100011, 8'b 01100111, 8'b 11100111, 8'b 11100110, 8'b 11000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00011000, 8'b 00011000, 8'b 11011011, 8'b 00111100, 8'b 11100111, 8'b 00111100, 8'b 11011011, 8'b 00011000, 8'b 00011000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 10000000, 8'b 11000000, 8'b 11100000, 8'b 11110000, 8'b 11111000, 8'b 11111110, 8'b 11111000, 8'b 11110000, 8'b 11100000, 8'b 11000000, 8'b 10000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000010, 8'b 00000110, 8'b 00001110, 8'b 00011110, 8'b 00111110, 8'b 11111110, 8'b 00111110, 8'b 00011110, 8'b 00001110, 8'b 00000110, 8'b 00000010, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00011000, 8'b 00111100, 8'b 01111110, 8'b 00011000, 8'b 00011000, 8'b 00011000, 8'b 01111110, 8'b 00111100, 8'b 00011000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 01100110, 8'b 01100110, 8'b 01100110, 8'b 01100110, 8'b 01100110, 8'b 01100110, 8'b 01100110, 8'b 00000000, 8'b 01100110, 8'b 01100110, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 01111111, 8'b 11011011, 8'b 11011011, 8'b 11011011, 8'b 01111011, 8'b 00011011, 8'b 00011011, 8'b 00011011, 8'b 00011011, 8'b 00011011, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 01111100, 8'b 11000110, 8'b 01100000, 8'b 00111000, 8'b 01101100, 8'b 11000110, 8'b 11000110, 8'b 01101100, 8'b 00111000, 8'b 00001100, 8'b 11000110, 8'b 01111100, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 11111110, 8'b 11111110, 8'b 11111110, 8'b 11111110, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00011000, 8'b 00111100, 8'b 01111110, 8'b 00011000, 8'b 00011000, 8'b 00011000, 8'b 01111110, 8'b 00111100, 8'b 00011000, 8'b 01111110, 8'b 00110000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00011000, 8'b 00111100, 8'b 01111110, 8'b 00011000, 8'b 00011000, 8'b 00011000, 8'b 00011000, 8'b 00011000, 8'b 00011000, 8'b 00011000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00011000, 8'b 00011000, 8'b 00011000, 8'b 00011000, 8'b 00011000, 8'b 00011000, 8'b 00011000, 8'b 01111110, 8'b 00111100, 8'b 00011000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00011000, 8'b 00001100, 8'b 11111110, 8'b 00001100, 8'b 00011000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00110000, 8'b 01100000, 8'b 11111110, 8'b 01100000, 8'b 00110000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 11000000, 8'b 11000000, 8'b 11000000, 8'b 11111110, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00100100, 8'b 01100110, 8'b 11111111, 8'b 01100110, 8'b 00100100, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00010000, 8'b 00111000, 8'b 00111000, 8'b 01111100, 8'b 01111100, 8'b 11111110, 8'b 11111110, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 11111110, 8'b 11111110, 8'b 01111100, 8'b 01111100, 8'b 00111000, 8'b 00111000, 8'b 00010000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00011000, 8'b 00111100, 8'b 00111100, 8'b 00111100, 8'b 00011000, 8'b 00011000, 8'b 00011000, 8'b 00000000, 8'b 00011000, 8'b 00011000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 01100110, 8'b 01100110, 8'b 01100110, 8'b 00100100, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 01101100, 8'b 01101100, 8'b 11111110, 8'b 01101100, 8'b 01101100, 8'b 01101100, 8'b 11111110, 8'b 01101100, 8'b 01101100, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00011000, 8'b 00011000, 8'b 01111100, 8'b 11000110, 8'b 11000010, 8'b 11000000, 8'b 01111100, 8'b 00000110, 8'b 00000110, 8'b 10000110, 8'b 11000110, 8'b 01111100, 8'b 00011000, 8'b 00011000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 11000010, 8'b 11000110, 8'b 00001100, 8'b 00011000, 8'b 00110000, 8'b 01100000, 8'b 11000110, 8'b 10000110, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00111000, 8'b 01101100, 8'b 01101100, 8'b 00111000, 8'b 01110110, 8'b 11011100, 8'b 11001100, 8'b 11001100, 8'b 11001100, 8'b 01110110, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00110000, 8'b 00110000, 8'b 00110000, 8'b 01100000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00001100, 8'b 00011000, 8'b 00110000, 8'b 00110000, 8'b 00110000, 8'b 00110000, 8'b 00110000, 8'b 00110000, 8'b 00011000, 8'b 00001100, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00110000, 8'b 00011000, 8'b 00001100, 8'b 00001100, 8'b 00001100, 8'b 00001100, 8'b 00001100, 8'b 00001100, 8'b 00011000, 8'b 00110000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 01100110, 8'b 00111100, 8'b 11111111, 8'b 00111100, 8'b 01100110, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00011000, 8'b 00011000, 8'b 01111110, 8'b 00011000, 8'b 00011000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00011000, 8'b 00011000, 8'b 00011000, 8'b 00110000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 01111110, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00011000, 8'b 00011000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000010, 8'b 00000110, 8'b 00001100, 8'b 00011000, 8'b 00110000, 8'b 01100000, 8'b 11000000, 8'b 10000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 01111100, 8'b 11000110, 8'b 11000110, 8'b 11001110, 8'b 11011110, 8'b 11110110, 8'b 11100110, 8'b 11000110, 8'b 11000110, 8'b 01111100, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00011000, 8'b 00111000, 8'b 01111000, 8'b 00011000, 8'b 00011000, 8'b 00011000, 8'b 00011000, 8'b 00011000, 8'b 00011000, 8'b 01111110, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 01111100, 8'b 11000110, 8'b 00000110, 8'b 00001100, 8'b 00011000, 8'b 00110000, 8'b 01100000, 8'b 11000000, 8'b 11000110, 8'b 11111110, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 01111100, 8'b 11000110, 8'b 00000110, 8'b 00000110, 8'b 00111100, 8'b 00000110, 8'b 00000110, 8'b 00000110, 8'b 11000110, 8'b 01111100, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00001100, 8'b 00011100, 8'b 00111100, 8'b 01101100, 8'b 11001100, 8'b 11111110, 8'b 00001100, 8'b 00001100, 8'b 00001100, 8'b 00011110, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 11111110, 8'b 11000000, 8'b 11000000, 8'b 11000000, 8'b 11111100, 8'b 00000110, 8'b 00000110, 8'b 00000110, 8'b 11000110, 8'b 01111100, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00111000, 8'b 01100000, 8'b 11000000, 8'b 11000000, 8'b 11111100, 8'b 11000110, 8'b 11000110, 8'b 11000110, 8'b 11000110, 8'b 01111100, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 11111110, 8'b 11000110, 8'b 00000110, 8'b 00000110, 8'b 00001100, 8'b 00011000, 8'b 00110000, 8'b 00110000, 8'b 00110000, 8'b 00110000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 01111100, 8'b 11000110, 8'b 11000110, 8'b 11000110, 8'b 01111100, 8'b 11000110, 8'b 11000110, 8'b 11000110, 8'b 11000110, 8'b 01111100, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 01111100, 8'b 11000110, 8'b 11000110, 8'b 11000110, 8'b 01111110, 8'b 00000110, 8'b 00000110, 8'b 00000110, 8'b 00001100, 8'b 01111000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00011000, 8'b 00011000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00011000, 8'b 00011000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00011000, 8'b 00011000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00011000, 8'b 00011000, 8'b 00110000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000110, 8'b 00001100, 8'b 00011000, 8'b 00110000, 8'b 01100000, 8'b 00110000, 8'b 00011000, 8'b 00001100, 8'b 00000110, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 01111110, 8'b 00000000, 8'b 00000000, 8'b 01111110, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 01100000, 8'b 00110000, 8'b 00011000, 8'b 00001100, 8'b 00000110, 8'b 00001100, 8'b 00011000, 8'b 00110000, 8'b 01100000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 01111100, 8'b 11000110, 8'b 11000110, 8'b 00001100, 8'b 00011000, 8'b 00011000, 8'b 00011000, 8'b 00000000, 8'b 00011000, 8'b 00011000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 01111100, 8'b 11000110, 8'b 11000110, 8'b 11000110, 8'b 11011110, 8'b 11011110, 8'b 11011110, 8'b 11011100, 8'b 11000000, 8'b 01111100, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00010000, 8'b 00111000, 8'b 01101100, 8'b 11000110, 8'b 11000110, 8'b 11111110, 8'b 11000110, 8'b 11000110, 8'b 11000110, 8'b 11000110, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 11111100, 8'b 01100110, 8'b 01100110, 8'b 01100110, 8'b 01111100, 8'b 01100110, 8'b 01100110, 8'b 01100110, 8'b 01100110, 8'b 11111100, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00111100, 8'b 01100110, 8'b 11000010, 8'b 11000000, 8'b 11000000, 8'b 11000000, 8'b 11000000, 8'b 11000010, 8'b 01100110, 8'b 00111100, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 11111000, 8'b 01101100, 8'b 01100110, 8'b 01100110, 8'b 01100110, 8'b 01100110, 8'b 01100110, 8'b 01100110, 8'b 01101100, 8'b 11111000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 11111110, 8'b 01100110, 8'b 01100010, 8'b 01101000, 8'b 01111000, 8'b 01101000, 8'b 01100000, 8'b 01100010, 8'b 01100110, 8'b 11111110, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 11111110, 8'b 01100110, 8'b 01100010, 8'b 01101000, 8'b 01111000, 8'b 01101000, 8'b 01100000, 8'b 01100000, 8'b 01100000, 8'b 11110000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00111100, 8'b 01100110, 8'b 11000010, 8'b 11000000, 8'b 11000000, 8'b 11011110, 8'b 11000110, 8'b 11000110, 8'b 01100110, 8'b 00111010, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 11000110, 8'b 11000110, 8'b 11000110, 8'b 11000110, 8'b 11111110, 8'b 11000110, 8'b 11000110, 8'b 11000110, 8'b 11000110, 8'b 11000110, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00111100, 8'b 00011000, 8'b 00011000, 8'b 00011000, 8'b 00011000, 8'b 00011000, 8'b 00011000, 8'b 00011000, 8'b 00011000, 8'b 00111100, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00011110, 8'b 00001100, 8'b 00001100, 8'b 00001100, 8'b 00001100, 8'b 00001100, 8'b 11001100, 8'b 11001100, 8'b 11001100, 8'b 01111000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 11100110, 8'b 01100110, 8'b 01100110, 8'b 01101100, 8'b 01111000, 8'b 01111000, 8'b 01101100, 8'b 01100110, 8'b 01100110, 8'b 11100110, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 11110000, 8'b 01100000, 8'b 01100000, 8'b 01100000, 8'b 01100000, 8'b 01100000, 8'b 01100000, 8'b 01100010, 8'b 01100110, 8'b 11111110, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 11000011, 8'b 11100111, 8'b 11111111, 8'b 11111111, 8'b 11011011, 8'b 11000011, 8'b 11000011, 8'b 11000011, 8'b 11000011, 8'b 11000011, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 11000110, 8'b 11100110, 8'b 11110110, 8'b 11111110, 8'b 11011110, 8'b 11001110, 8'b 11000110, 8'b 11000110, 8'b 11000110, 8'b 11000110, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 01111100, 8'b 11000110, 8'b 11000110, 8'b 11000110, 8'b 11000110, 8'b 11000110, 8'b 11000110, 8'b 11000110, 8'b 11000110, 8'b 01111100, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 11111100, 8'b 01100110, 8'b 01100110, 8'b 01100110, 8'b 01111100, 8'b 01100000, 8'b 01100000, 8'b 01100000, 8'b 01100000, 8'b 11110000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 01111100, 8'b 11000110, 8'b 11000110, 8'b 11000110, 8'b 11000110, 8'b 11000110, 8'b 11000110, 8'b 11010110, 8'b 11011110, 8'b 01111100, 8'b 00001100, 8'b 00001110, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 11111100, 8'b 01100110, 8'b 01100110, 8'b 01100110, 8'b 01111100, 8'b 01101100, 8'b 01100110, 8'b 01100110, 8'b 01100110, 8'b 11100110, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 01111100, 8'b 11000110, 8'b 11000110, 8'b 01100000, 8'b 00111000, 8'b 00001100, 8'b 00000110, 8'b 11000110, 8'b 11000110, 8'b 01111100, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 11111111, 8'b 11011011, 8'b 10011001, 8'b 00011000, 8'b 00011000, 8'b 00011000, 8'b 00011000, 8'b 00011000, 8'b 00011000, 8'b 00111100, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 11000110, 8'b 11000110, 8'b 11000110, 8'b 11000110, 8'b 11000110, 8'b 11000110, 8'b 11000110, 8'b 11000110, 8'b 11000110, 8'b 01111100, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 11000011, 8'b 11000011, 8'b 11000011, 8'b 11000011, 8'b 11000011, 8'b 11000011, 8'b 11000011, 8'b 01100110, 8'b 00111100, 8'b 00011000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 11000011, 8'b 11000011, 8'b 11000011, 8'b 11000011, 8'b 11000011, 8'b 11011011, 8'b 11011011, 8'b 11111111, 8'b 01100110, 8'b 01100110, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 11000011, 8'b 11000011, 8'b 01100110, 8'b 00111100, 8'b 00011000, 8'b 00011000, 8'b 00111100, 8'b 01100110, 8'b 11000011, 8'b 11000011, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 11000011, 8'b 11000011, 8'b 11000011, 8'b 01100110, 8'b 00111100, 8'b 00011000, 8'b 00011000, 8'b 00011000, 8'b 00011000, 8'b 00111100, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 11111111, 8'b 11000011, 8'b 10000110, 8'b 00001100, 8'b 00011000, 8'b 00110000, 8'b 01100000, 8'b 11000001, 8'b 11000011, 8'b 11111111, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00111100, 8'b 00110000, 8'b 00110000, 8'b 00110000, 8'b 00110000, 8'b 00110000, 8'b 00110000, 8'b 00110000, 8'b 00110000, 8'b 00111100, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 10000000, 8'b 11000000, 8'b 11100000, 8'b 01110000, 8'b 00111000, 8'b 00011100, 8'b 00001110, 8'b 00000110, 8'b 00000010, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00111100, 8'b 00001100, 8'b 00001100, 8'b 00001100, 8'b 00001100, 8'b 00001100, 8'b 00001100, 8'b 00001100, 8'b 00001100, 8'b 00111100, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00010000, 8'b 00111000, 8'b 01101100, 8'b 11000110, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 11111111, 8'b 00000000, 8'b 00000000, 8'b 00110000, 8'b 00110000, 8'b 00011000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 01111000, 8'b 00001100, 8'b 01111100, 8'b 11001100, 8'b 11001100, 8'b 11001100, 8'b 01110110, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 11100000, 8'b 01100000, 8'b 01100000, 8'b 01111000, 8'b 01101100, 8'b 01100110, 8'b 01100110, 8'b 01100110, 8'b 01100110, 8'b 01111100, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 01111100, 8'b 11000110, 8'b 11000000, 8'b 11000000, 8'b 11000000, 8'b 11000110, 8'b 01111100, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00011100, 8'b 00001100, 8'b 00001100, 8'b 00111100, 8'b 01101100, 8'b 11001100, 8'b 11001100, 8'b 11001100, 8'b 11001100, 8'b 01110110, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 01111100, 8'b 11000110, 8'b 11111110, 8'b 11000000, 8'b 11000000, 8'b 11000110, 8'b 01111100, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00111000, 8'b 01101100, 8'b 01100100, 8'b 01100000, 8'b 11110000, 8'b 01100000, 8'b 01100000, 8'b 01100000, 8'b 01100000, 8'b 11110000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 01110110, 8'b 11001100, 8'b 11001100, 8'b 11001100, 8'b 11001100, 8'b 11001100, 8'b 01111100, 8'b 00001100, 8'b 11001100, 8'b 01111000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 11100000, 8'b 01100000, 8'b 01100000, 8'b 01101100, 8'b 01110110, 8'b 01100110, 8'b 01100110, 8'b 01100110, 8'b 01100110, 8'b 11100110, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00011000, 8'b 00011000, 8'b 00000000, 8'b 00111000, 8'b 00011000, 8'b 00011000, 8'b 00011000, 8'b 00011000, 8'b 00011000, 8'b 00111100, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000110, 8'b 00000110, 8'b 00000000, 8'b 00001110, 8'b 00000110, 8'b 00000110, 8'b 00000110, 8'b 00000110, 8'b 00000110, 8'b 00000110, 8'b 01100110, 8'b 01100110, 8'b 00111100, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 11100000, 8'b 01100000, 8'b 01100000, 8'b 01100110, 8'b 01101100, 8'b 01111000, 8'b 01111000, 8'b 01101100, 8'b 01100110, 8'b 11100110, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00111000, 8'b 00011000, 8'b 00011000, 8'b 00011000, 8'b 00011000, 8'b 00011000, 8'b 00011000, 8'b 00011000, 8'b 00011000, 8'b 00111100, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 11100110, 8'b 11111111, 8'b 11011011, 8'b 11011011, 8'b 11011011, 8'b 11011011, 8'b 11011011, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 11011100, 8'b 01100110, 8'b 01100110, 8'b 01100110, 8'b 01100110, 8'b 01100110, 8'b 01100110, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 01111100, 8'b 11000110, 8'b 11000110, 8'b 11000110, 8'b 11000110, 8'b 11000110, 8'b 01111100, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 11011100, 8'b 01100110, 8'b 01100110, 8'b 01100110, 8'b 01100110, 8'b 01100110, 8'b 01111100, 8'b 01100000, 8'b 01100000, 8'b 11110000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 01110110, 8'b 11001100, 8'b 11001100, 8'b 11001100, 8'b 11001100, 8'b 11001100, 8'b 01111100, 8'b 00001100, 8'b 00001100, 8'b 00011110, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 11011100, 8'b 01110110, 8'b 01100110, 8'b 01100000, 8'b 01100000, 8'b 01100000, 8'b 11110000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 01111100, 8'b 11000110, 8'b 01100000, 8'b 00111000, 8'b 00001100, 8'b 11000110, 8'b 01111100, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00010000, 8'b 00110000, 8'b 00110000, 8'b 11111100, 8'b 00110000, 8'b 00110000, 8'b 00110000, 8'b 00110000, 8'b 00110110, 8'b 00011100, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 11001100, 8'b 11001100, 8'b 11001100, 8'b 11001100, 8'b 11001100, 8'b 11001100, 8'b 01110110, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 11000011, 8'b 11000011, 8'b 11000011, 8'b 11000011, 8'b 01100110, 8'b 00111100, 8'b 00011000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 11000011, 8'b 11000011, 8'b 11000011, 8'b 11011011, 8'b 11011011, 8'b 11111111, 8'b 01100110, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 11000011, 8'b 01100110, 8'b 00111100, 8'b 00011000, 8'b 00111100, 8'b 01100110, 8'b 11000011, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 11000110, 8'b 11000110, 8'b 11000110, 8'b 11000110, 8'b 11000110, 8'b 11000110, 8'b 01111110, 8'b 00000110, 8'b 00001100, 8'b 11111000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 11111110, 8'b 11001100, 8'b 00011000, 8'b 00110000, 8'b 01100000, 8'b 11000110, 8'b 11111110, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00001110, 8'b 00011000, 8'b 00011000, 8'b 00011000, 8'b 01110000, 8'b 00011000, 8'b 00011000, 8'b 00011000, 8'b 00011000, 8'b 00001110, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00011000, 8'b 00011000, 8'b 00011000, 8'b 00011000, 8'b 00000000, 8'b 00011000, 8'b 00011000, 8'b 00011000, 8'b 00011000, 8'b 00011000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 01110000, 8'b 00011000, 8'b 00011000, 8'b 00011000, 8'b 00001110, 8'b 00011000, 8'b 00011000, 8'b 00011000, 8'b 00011000, 8'b 01110000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 01110110, 8'b 11011100, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00010000, 8'b 00111000, 8'b 01101100, 8'b 11000110, 8'b 11000110, 8'b 11000110, 8'b 11111110, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000, 8'b 00000000}; 

//  2^11-by-8
//  0
//  1
//  2
//  3
//  4
//  5
//  6
//  7
//  8
//  9
//  a
//  b
//  c
//  d
//  e
//  f
//  code x01
//  0
//  1
//  2  ******
//  3 *      *
//  4 * *  * *
//  5 *      *
//  6 *      *
//  7 * **** *
//  8 *  **  *
//  9 *      *
//  a *      *
//  b  ******
//  c
//  d
//  e
//  f
//  code x02
//  0
//  1
//  2  ******
//  3 ********
//  4 ** ** **
//  5 ********
//  6 ********
//  7 **    **
//  8 ***  ***
//  9 ********
//  a ********
//  b  ******
//  c
//  d
//  e
//  f
//  code x03
//  0
//  1
//  2
//  3
//  4  ** **
//  5 *******
//  6 *******
//  7 *******
//  8 *******
//  9  *****
//  a   ***
//  b    *
//  c
//  d
//  e
//  f
//  code x04
//  0
//  1
//  2
//  3
//  4    *
//  5   ***
//  6  *****
//  7 *******
//  8  *****
//  9   ***
//  a    *
//  b
//  c
//  d
//  e
//  f
//  code x05
//  0
//  1
//  2
//  3    **
//  4   ****
//  5   ****
//  6 ***  ***
//  7 ***  ***
//  8 ***  ***
//  9    **
//  a    **
//  b   ****
//  c
//  d
//  e
//  f
//  code x06
//  0
//  1
//  2
//  3    **
//  4   ****
//  5  ******
//  6 ********
//  7 ********
//  8  ******
//  9    **
//  a    **
//  b   ****
//  c
//  d
//  e
//  f
//  code x07
//  0
//  1
//  2
//  3
//  4
//  5
//  6    **
//  7   ****
//  8   ****
//  9    **
//  a
//  b
//  c
//  d
//  e
//  f
//  code x08
//  0 ********
//  1 ********
//  2 ********
//  3 ********
//  4 ********
//  5 ********
//  6 ***  ***
//  7 **    **
//  8 **    **
//  9 ***  ***
//  a ********
//  b ********
//  c ********
//  d ********
//  e ********
//  f ********
//  code x09
//  0
//  1
//  2
//  3
//  4
//  5   ****
//  6  **  **
//  7  *    *
//  8  *    *
//  9  **  **
//  a   ****
//  b
//  c
//  d
//  e
//  f
//  code x0a
//  0 ********
//  1 ********
//  2 ********
//  3 ********
//  4 ********
//  5 **    **
//  6 *  **  *
//  7 * **** *
//  8 * **** *
//  9 *  **  *
//  a **    **
//  b ********
//  c ********
//  d ********
//  e ********
//  f ********
//  code x0b
//  0
//  1
//  2    ****
//  3     ***
//  4    ** *
//  5   **  *
//  6  ****
//  7 **  **
//  8 **  **
//  9 **  **
//  a **  **
//  b  ****
//  c
//  d
//  e
//  f
//  code x0c
//  0
//  1
//  2   ****
//  3  **  **
//  4  **  **
//  5  **  **
//  6  **  **
//  7   ****
//  8    **
//  9  ******
//  a    **
//  b    **
//  c
//  d
//  e
//  f
//  code x0d
//  0
//  1
//  2   ******
//  3   **  **
//  4   ******
//  5   **
//  6   **
//  7   **
//  8   **
//  9  ***
//  a ****
//  b ***
//  c
//  d
//  e
//  f
//  code x0e
//  0
//  1
//  2  *******
//  3  **   **
//  4  *******
//  5  **   **
//  6  **   **
//  7  **   **
//  8  **   **
//  9  **  ***
//  a ***  ***
//  b ***  **
//  c **
//  d
//  e
//  f
//  code x0f
//  0
//  1
//  2
//  3    **
//  4    **
//  5 ** ** **
//  6   ****
//  7 ***  ***
//  8   ****
//  9 ** ** **
//  a    **
//  b    **
//  c
//  d
//  e
//  f
//  code x10
//  0
//  1 *
//  2 **
//  3 ***
//  4 ****
//  5 *****
//  6 *******
//  7 *****
//  8 ****
//  9 ***
//  a **
//  b *
//  c
//  d
//  e
//  f
//  code x11
//  0
//  1       *
//  2      **
//  3     ***
//  4    ****
//  5   *****
//  6 *******
//  7   *****
//  8    ****
//  9     ***
//  a      **
//  b       *
//  c
//  d
//  e
//  f
//  code x12
//  0
//  1
//  2    **
//  3   ****
//  4  ******
//  5    **
//  6    **
//  7    **
//  8  ******
//  9   ****
//  a    **
//  b
//  c
//  d
//  e
//  f
//  code x13
//  0
//  1
//  2  **  **
//  3  **  **
//  4  **  **
//  5  **  **
//  6  **  **
//  7  **  **
//  8  **  **
//  9
//  a  **  **
//  b  **  **
//  c
//  d
//  e
//  f
//  code x14
//  0
//  1
//  2  *******
//  3 ** ** **
//  4 ** ** **
//  5 ** ** **
//  6  **** **
//  7    ** **
//  8    ** **
//  9    ** **
//  a    ** **
//  b    ** **
//  c
//  d
//  e
//  f
//  code x15
//  0
//  1  *****
//  2 **   **
//  3  **
//  4   ***
//  5  ** **
//  6 **   **
//  7 **   **
//  8  ** **
//  9   ***
//  a     **
//  b **   **
//  c  *****
//  d
//  e
//  f
//  code x16
//  0
//  1
//  2
//  3
//  4
//  5
//  6
//  7
//  8 *******
//  9 *******
//  a *******
//  b *******
//  c
//  d
//  e
//  f
//  code x17
//  0
//  1
//  2    **
//  3   ****
//  4  ******
//  5    **
//  6    **
//  7    **
//  8  ******
//  9   ****
//  a    **
//  b  ******
//  c
//  d
//  e
//  f
//  code x18
//  0
//  1
//  2    **
//  3   ****
//  4  ******
//  5    **
//  6    **
//  7    **
//  8    **
//  9    **
//  a    **
//  b    **
//  c
//  d
//  e
//  f
//  code x19
//  0
//  1
//  2    **
//  3    **
//  4    **
//  5    **
//  6    **
//  7    **
//  8    **
//  9  ******
//  a   ****
//  b    **
//  c
//  d
//  e
//  f
//  code x1a
//  0
//  1
//  2
//  3
//  4
//  5    **
//  6     **
//  7 *******
//  8     **
//  9    **
//  a
//  b
//  c
//  d
//  e
//  f
//  code x1b
//  0
//  1
//  2
//  3
//  4
//  5   **
//  6  **
//  7 *******
//  8  **
//  9   **
//  a
//  b
//  c
//  d
//  e
//  f
//  code x1c
//  0
//  1
//  2
//  3
//  4
//  5
//  6 **
//  7 **
//  8 **
//  9 *******
//  a
//  b
//  c
//  d
//  e
//  f
//  code x1d
//  0
//  1
//  2
//  3
//  4
//  5   *  *
//  6  **  **
//  7 ********
//  8  **  **
//  9   *  *
//  a
//  b
//  c
//  d
//  e
//  f
//  code x1e
//  0
//  1
//  2
//  3
//  4    *
//  5   ***
//  6   ***
//  7  *****
//  8  *****
//  9 *******
//  a *******
//  b
//  c
//  d
//  e
//  f
//  code x1f
//  0
//  1
//  2
//  3
//  4 *******
//  5 *******
//  6  *****
//  7  *****
//  8   ***
//  9   ***
//  a    *
//  b
//  c
//  d
//  e
//  f
//  code x20
//  0
//  1
//  2
//  3
//  4
//  5
//  6
//  7
//  8
//  9
//  a
//  b
//  c
//  d
//  e
//  f
//  code x21
//  0
//  1
//  2    **
//  3   ****
//  4   ****
//  5   ****
//  6    **
//  7    **
//  8    **
//  9
//  a    **
//  b    **
//  c
//  d
//  e
//  f
//  code x22
//  0
//  1  **  **
//  2  **  **
//  3  **  **
//  4   *  *
//  5
//  6
//  7
//  8
//  9
//  a
//  b
//  c
//  d
//  e
//  f
//  code x23
//  0
//  1
//  2
//  3  ** **
//  4  ** **
//  5 *******
//  6  ** **
//  7  ** **
//  8  ** **
//  9 *******
//  a  ** **
//  b  ** **
//  c
//  d
//  e
//  f
//  code x24
//  0     **
//  1     **
//  2   *****
//  3  **   **
//  4  **    *
//  5  **
//  6   *****
//  7       **
//  8       **
//  9  *    **
//  a  **   **
//  b   *****
//  c     **
//  d     **
//  e
//  f
//  code x25
//  0
//  1
//  2
//  3
//  4 **    *
//  5 **   **
//  6     **
//  7    **
//  8   **
//  9  **
//  a **   **
//  b *    **
//  c
//  d
//  e
//  f
//  code x26
//  0
//  1
//  2   ***
//  3  ** **
//  4  ** **
//  5   ***
//  6  *** **
//  7 ** ***
//  8 **  **
//  9 **  **
//  a **  **
//  b  *** **
//  c
//  d
//  e
//  f
//  code x27
//  0
//  1   **
//  2   **
//  3   **
//  4  **
//  5
//  6
//  7
//  8
//  9
//  a
//  b
//  c
//  d
//  e
//  f
//  code x28
//  0
//  1
//  2     **
//  3    **
//  4   **
//  5   **
//  6   **
//  7   **
//  8   **
//  9   **
//  a    **
//  b     **
//  c
//  d
//  e
//  f
//  code x29
//  0
//  1
//  2   **
//  3    **
//  4     **
//  5     **
//  6     **
//  7     **
//  8     **
//  9     **
//  a    **
//  b   **
//  c
//  d
//  e
//  f
//  code x2a
//  0
//  1
//  2
//  3
//  4
//  5  **  **
//  6   ****
//  7 ********
//  8   ****
//  9  **  **
//  a
//  b
//  c
//  d
//  e
//  f
//  code x2b
//  0
//  1
//  2
//  3
//  4
//  5    **
//  6    **
//  7  ******
//  8    **
//  9    **
//  a
//  b
//  c
//  d
//  e
//  f
//  code x2c
//  0
//  1
//  2
//  3
//  4
//  5
//  6
//  7
//  8
//  9    **
//  a    **
//  b    **
//  c   **
//  d
//  e
//  f
//  code x2d
//  0
//  1
//  2
//  3
//  4
//  5
//  6
//  7  ******
//  8
//  9
//  a
//  b
//  c
//  d
//  e
//  f
//  code x2e
//  0
//  1
//  2
//  3
//  4
//  5
//  6
//  7
//  8
//  9
//  a    **
//  b    **
//  c
//  d
//  e
//  f
//  code x2f
//  0
//  1
//  2
//  3
//  4       *
//  5      **
//  6     **
//  7    **
//  8   **
//  9  **
//  a **
//  b *
//  c
//  d
//  e
//  f
//  code x30
//  0
//  1
//  2  *****
//  3 **   **
//  4 **   **
//  5 **  ***
//  6 ** ****
//  7 **** **
//  8 ***  **
//  9 **   **
//  a **   **
//  b  *****
//  c
//  d
//  e
//  f
//  code x31
//  0
//  1
//  2
//  3
//  4    **
//  5   ***
//  6  ****
//  7    **
//  8    **
//  9    **
//  a    **
//  b    **
//  c    **
//  d  ******
//  e
//  f
//  code x32
//  0
//  1
//  2  *****
//  3 **   **
//  4      **
//  5     **
//  6    **
//  7   **
//  8  **
//  9 **
//  a **   **
//  b *******
//  c
//  d
//  e
//  f
//  code x33
//  0
//  1
//  2  *****
//  3 **   **
//  4      **
//  5      **
//  6   ****
//  7      **
//  8      **
//  9      **
//  a **   **
//  b  *****
//  c
//  d
//  e
//  f
//  code x34
//  0
//  1
//  2     **
//  3    ***
//  4   ****
//  5  ** **
//  6 **  **
//  7 *******
//  8     **
//  9     **
//  a     **
//  b    ****
//  c
//  d
//  e
//  f
//  code x35
//  0
//  1
//  2 *******
//  3 **
//  4 **
//  5 **
//  6 ******
//  7      **
//  8      **
//  9      **
//  a **   **
//  b  *****
//  c
//  d
//  e
//  f
//  code x36
//  0
//  1
//  2   ***
//  3  **
//  4 **
//  5 **
//  6 ******
//  7 **   **
//  8 **   **
//  9 **   **
//  a **   **
//  b  *****
//  c
//  d
//  e
//  f
//  code x37
//  0
//  1
//  2 *******
//  3 **   **
//  4      **
//  5      **
//  6     **
//  7    **
//  8   **
//  9   **
//  a   **
//  b   **
//  c
//  d
//  e
//  f
//  code x38
//  0
//  1
//  2  *****
//  3 **   **
//  4 **   **
//  5 **   **
//  6  *****
//  7 **   **
//  8 **   **
//  9 **   **
//  a **   **
//  b  *****
//  c
//  d
//  e
//  f
//  code x39
//  0
//  1
//  2  *****
//  3 **   **
//  4 **   **
//  5 **   **
//  6  ******
//  7      **
//  8      **
//  9      **
//  a     **
//  b  ****
//  c
//  d
//  e
//  f
//  code x3a
//  0
//  1
//  2
//  3
//  4    **
//  5    **
//  6
//  7
//  8
//  9    **
//  a    **
//  b
//  c
//  d
//  e
//  f
//  code x3b
//  0
//  1
//  2
//  3
//  4    **
//  5    **
//  6
//  7
//  8
//  9    **
//  a    **
//  b   **
//  c
//  d
//  e
//  f
//  code x3c
//  0
//  1
//  2
//  3      **
//  4     **
//  5    **
//  6   **
//  7  **
//  8   **
//  9    **
//  a     **
//  b      **
//  c
//  d
//  e
//  f
//  code x3d
//  0
//  1
//  2
//  3
//  4
//  5  ******
//  6
//  7
//  8  ******
//  9
//  a
//  b
//  c
//  d
//  e
//  f
//  code x3e
//  0
//  1
//  2
//  3  **
//  4   **
//  5    **
//  6     **
//  7      **
//  8     **
//  9    **
//  a   **
//  b  **
//  c
//  d
//  e
//  f
//  code x3f
//  0
//  1
//  2  *****
//  3 **   **
//  4 **   **
//  5     **
//  6    **
//  7    **
//  8    **
//  9
//  a    **
//  b    **
//  c
//  d
//  e
//  f
//  code x40
//  0
//  1
//  2  *****
//  3 **   **
//  4 **   **
//  5 **   **
//  6 ** ****
//  7 ** ****
//  8 ** ****
//  9 ** ***
//  a **
//  b  *****
//  c
//  d
//  e
//  f
//  code x41
//  0
//  1
//  2    *
//  3   ***
//  4  ** **
//  5 **   **
//  6 **   **
//  7 *******
//  8 **   **
//  9 **   **
//  a **   **
//  b **   **
//  c
//  d
//  e
//  f
//  code x42
//  0
//  1
//  2 ******
//  3  **  **
//  4  **  **
//  5  **  **
//  6  *****
//  7  **  **
//  8  **  **
//  9  **  **
//  a  **  **
//  b ******
//  c
//  d
//  e
//  f
//  code x43
//  0
//  1
//  2   ****
//  3  **  **
//  4 **    *
//  5 **
//  6 **
//  7 **
//  8 **
//  9 **    *
//  a  **  **
//  b   ****
//  c
//  d
//  e
//  f
//  code x44
//  0
//  1
//  2 *****
//  3  ** **
//  4  **  **
//  5  **  **
//  6  **  **
//  7  **  **
//  8  **  **
//  9  **  **
//  a  ** **
//  b *****
//  c
//  d
//  e
//  f
//  code x45
//  0
//  1
//  2 *******
//  3  **  **
//  4  **   *
//  5  ** *
//  6  ****
//  7  ** *
//  8  **
//  9  **   *
//  a  **  **
//  b *******
//  c
//  d
//  e
//  f
//  code x46
//  0
//  1
//  2 *******
//  3  **  **
//  4  **   *
//  5  ** *
//  6  ****
//  7  ** *
//  8  **
//  9  **
//  a  **
//  b ****
//  c
//  d
//  e
//  f
//  code x47
//  0
//  1
//  2   ****
//  3  **  **
//  4 **    *
//  5 **
//  6 **
//  7 ** ****
//  8 **   **
//  9 **   **
//  a  **  **
//  b   *** *
//  c
//  d
//  e
//  f
//  code x48
//  0
//  1
//  2 **   **
//  3 **   **
//  4 **   **
//  5 **   **
//  6 *******
//  7 **   **
//  8 **   **
//  9 **   **
//  a **   **
//  b **   **
//  c
//  d
//  e
//  f
//  code x49
//  0
//  1
//  2   ****
//  3    **
//  4    **
//  5    **
//  6    **
//  7    **
//  8    **
//  9    **
//  a    **
//  b   ****
//  c
//  d
//  e
//  f
//  code x4a
//  0
//  1
//  2    ****
//  3     **
//  4     **
//  5     **
//  6     **
//  7     **
//  8 **  **
//  9 **  **
//  a **  **
//  b  ****
//  c
//  d
//  e
//  f
//  code x4b
//  0
//  1
//  2 ***  **
//  3  **  **
//  4  **  **
//  5  ** **
//  6  ****
//  7  ****
//  8  ** **
//  9  **  **
//  a  **  **
//  b ***  **
//  c
//  d
//  e
//  f
//  code x4c
//  0
//  1
//  2 ****
//  3  **
//  4  **
//  5  **
//  6  **
//  7  **
//  8  **
//  9  **   *
//  a  **  **
//  b *******
//  c
//  d
//  e
//  f
//  code x4d
//  0
//  1
//  2 **    **
//  3 ***  ***
//  4 ********
//  5 ********
//  6 ** ** **
//  7 **    **
//  8 **    **
//  9 **    **
//  a **    **
//  b **    **
//  c
//  d
//  e
//  f
//  code x4e
//  0
//  1
//  2 **   **
//  3 ***  **
//  4 **** **
//  5 *******
//  6 ** ****
//  7 **  ***
//  8 **   **
//  9 **   **
//  a **   **
//  b **   **
//  c
//  d
//  e
//  f
//  code x4f
//  0
//  1
//  2  *****
//  3 **   **
//  4 **   **
//  5 **   **
//  6 **   **
//  7 **   **
//  8 **   **
//  9 **   **
//  a **   **
//  b  *****
//  c
//  d
//  e
//  f
//  code x50
//  0
//  1
//  2 ******
//  3  **  **
//  4  **  **
//  5  **  **
//  6  *****
//  7  **
//  8  **
//  9  **
//  a  **
//  b ****
//  c
//  d
//  e
//  f
//  code x510
//  0
//  1
//  2  *****
//  3 **   **
//  4 **   **
//  5 **   **
//  6 **   **
//  7 **   **
//  8 **   **
//  9 ** * **
//  a ** ****
//  b  *****
//  c     **
//  d     ***
//  e
//  f
//  code x52
//  0
//  1
//  2 ******
//  3  **  **
//  4  **  **
//  5  **  **
//  6  *****
//  7  ** **
//  8  **  **
//  9  **  **
//  a  **  **
//  b ***  **
//  c
//  d
//  e
//  f
//  code x53
//  0
//  1
//  2  *****
//  3 **   **
//  4 **   **
//  5  **
//  6   ***
//  7     **
//  8      **
//  9 **   **
//  a **   **
//  b  *****
//  c
//  d
//  e
//  f
//  code x54
//  0
//  1
//  2 ********
//  3 ** ** **
//  4 *  **  *
//  5    **
//  6    **
//  7    **
//  8    **
//  9    **
//  a    **
//  b   ****
//  c
//  d
//  e
//  f
//  code x55
//  0
//  1
//  2 **   **
//  3 **   **
//  4 **   **
//  5 **   **
//  6 **   **
//  7 **   **
//  8 **   **
//  9 **   **
//  a **   **
//  b  *****
//  c
//  d
//  e
//  f
//  code x56
//  0
//  1
//  2 **    **
//  3 **    **
//  4 **    **
//  5 **    **
//  6 **    **
//  7 **    **
//  8 **    **
//  9  **  **
//  a   ****
//  b    **
//  c
//  d
//  e
//  f
//  code x57
//  0
//  1
//  2 **    **
//  3 **    **
//  4 **    **
//  5 **    **
//  6 **    **
//  7 ** ** **
//  8 ** ** **
//  9 ********
//  a  **  **
//  b  **  **
//  c
//  d
//  e
//  f
//  code x58
//  0
//  1
//  2 **    **
//  3 **    **
//  4  **  **
//  5   ****
//  6    **
//  7    **
//  8   ****
//  9  **  **
//  a **    **
//  b **    **
//  c
//  d
//  e
//  f
//  code x59
//  0
//  1
//  2 **    **
//  3 **    **
//  4 **    **
//  5  **  **
//  6   ****
//  7    **
//  8    **
//  9    **
//  a    **
//  b   ****
//  c
//  d
//  e
//  f
//  code x5a
//  0
//  1
//  2 ********
//  3 **    **
//  4 *    **
//  5     **
//  6    **
//  7   **
//  8  **
//  9 **     *
//  a **    **
//  b ********
//  c
//  d
//  e
//  f
//  code x5b
//  0
//  1
//  2   ****
//  3   **
//  4   **
//  5   **
//  6   **
//  7   **
//  8   **
//  9   **
//  a   **
//  b   ****
//  c
//  d
//  e
//  f
//  code x5c
//  0
//  1
//  2
//  3 *
//  4 **
//  5 ***
//  6  ***
//  7   ***
//  8    ***
//  9     ***
//  a      **
//  b       *
//  c
//  d
//  e
//  f
//  code x5d
//  0
//  1
//  2   ****
//  3     **
//  4     **
//  5     **
//  6     **
//  7     **
//  8     **
//  9     **
//  a     **
//  b   ****
//  c
//  d
//  e
//  f
//  code x5e
//  0    *
//  1   ***
//  2  ** **
//  3 **   **
//  4
//  5
//  6
//  7
//  8
//  9
//  a
//  b
//  c
//  d
//  e
//  f
//  code x5f
//  0
//  1
//  2
//  3
//  4
//  5
//  6
//  7
//  8
//  9
//  a
//  b
//  c
//  d ********
//  e
//  f
//  code x60
//  0   **
//  1   **
//  2    **
//  3
//  4
//  5
//  6
//  7
//  8
//  9
//  a
//  b
//  c
//  d
//  e
//  f
//  code x61
//  0
//  1
//  2
//  3
//  4
//  5  ****
//  6     **
//  7  *****
//  8 **  **
//  9 **  **
//  a **  **
//  b  *** **
//  c
//  d
//  e
//  f
//  code x62
//  0
//  1
//  2  ***
//  3   **
//  4   **
//  5   ****
//  6   ** **
//  7   **  **
//  8   **  **
//  9   **  **
//  a   **  **
//  b   *****
//  c
//  d
//  e
//  f
//  code x63
//  0
//  1
//  2
//  3
//  4
//  5  *****
//  6 **   **
//  7 **
//  8 **
//  9 **
//  a **   **
//  b  *****
//  c
//  d
//  e
//  f
//  code x64
//  0
//  1
//  2    ***
//  3     **
//  4     **
//  5   ****
//  6  ** **
//  7 **  **
//  8 **  **
//  9 **  **
//  a **  **
//  b  *** **
//  c
//  d
//  e
//  f
//  code x65
//  0
//  1
//  2
//  3
//  4
//  5  *****
//  6 **   **
//  7 *******
//  8 **
//  9 **
//  a **   **
//  b  *****
//  c
//  d
//  e
//  f
//  code x66
//  0
//  1
//  2   ***
//  3  ** **
//  4  **  *
//  5  **
//  6 ****
//  7  **
//  8  **
//  9  **
//  a  **
//  b ****
//  c
//  d
//  e
//  f
//  code x67
//  0
//  1
//  2
//  3
//  4
//  5  *** **
//  6 **  **
//  7 **  **
//  8 **  **
//  9 **  **
//  a **  **
//  b  *****
//  c     **
//  d **  **
//  e  ****
//  f
//  code x68
//  0
//  1
//  2 ***
//  3  **
//  4  **
//  5  ** **
//  6  *** **
//  7  **  **
//  8  **  **
//  9  **  **
//  a  **  **
//  b ***  **
//  c
//  d
//  e
//  f
//  code x69
//  0
//  1
//  2    **
//  3    **
//  4
//  5   ***
//  6    **
//  7    **
//  8    **
//  9    **
//  a    **
//  b   ****
//  c
//  d
//  e
//  f
//  code x6a
//  0
//  1
//  2      **
//  3      **
//  4
//  5     ***
//  6      **
//  7      **
//  8      **
//  9      **
//  a      **
//  b      **
//  c  **  **
//  d  **  **
//  e   ****
//  f
//  code x6b
//  0
//  1
//  2 ***
//  3  **
//  4  **
//  5  **  **
//  6  ** **
//  7  ****
//  8  ****
//  9  ** **
//  a  **  **
//  b ***  **
//  c
//  d
//  e
//  f
//  code x6c
//  0
//  1
//  2   ***
//  3    **
//  4    **
//  5    **
//  6    **
//  7    **
//  8    **
//  9    **
//  a    **
//  b   ****
//  c
//  d
//  e
//  f
//  code x6d
//  0
//  1
//  2
//  3
//  4
//  5 ***  **
//  6 ********
//  7 ** ** **
//  8 ** ** **
//  9 ** ** **
//  a ** ** **
//  b ** ** **
//  c
//  d
//  e
//  f
//  code x6e
//  0
//  1
//  2
//  3
//  4
//  5 ** ***
//  6  **  **
//  7  **  **
//  8  **  **
//  9  **  **
//  a  **  **
//  b  **  **
//  c
//  d
//  e
//  f
//  code x6f
//  0
//  1
//  2
//  3
//  4
//  5  *****
//  6 **   **
//  7 **   **
//  8 **   **
//  9 **   **
//  a **   **
//  b  *****
//  c
//  d
//  e
//  f
//  code x70
//  0
//  1
//  2
//  3
//  4
//  5 ** ***
//  6  **  **
//  7  **  **
//  8  **  **
//  9  **  **
//  a  **  **
//  b  *****
//  c  **
//  d  **
//  e ****
//  f
//  code x71
//  0
//  1
//  2
//  3
//  4
//  5  *** **
//  6 **  **
//  7 **  **
//  8 **  **
//  9 **  **
//  a **  **
//  b  *****
//  c     **
//  d     **
//  e    ****
//  f
//  code x72
//  0
//  1
//  2
//  3
//  4
//  5 ** ***
//  6  *** **
//  7  **  **
//  8  **
//  9  **
//  a  **
//  b ****
//  c
//  d
//  e
//  f
//  code x73
//  0
//  1
//  2
//  3
//  4
//  5  *****
//  6 **   **
//  7  **
//  8   ***
//  9     **
//  a **   **
//  b  *****
//  c
//  d
//  e
//  f
//  code x74
//  0
//  1
//  2    *
//  3   **
//  4   **
//  5 ******
//  6   **
//  7   **
//  8   **
//  9   **
//  a   ** **
//  b    ***
//  c
//  d
//  e
//  f
//  code x75
//  0
//  1
//  2
//  3
//  4
//  5 **  **
//  6 **  **
//  7 **  **
//  8 **  **
//  9 **  **
//  a **  **
//  b  *** **
//  c
//  d
//  e
//  f
//  code x76
//  0
//  1
//  2
//  3
//  4
//  5 **    **
//  6 **    **
//  7 **    **
//  8 **    **
//  9  **  **
//  a   ****
//  b    **
//  c
//  d
//  e
//  f
//  code x77
//  0
//  1
//  2
//  3
//  4
//  5 **    **
//  6 **    **
//  7 **    **
//  8 ** ** **
//  9 ** ** **
//  a ********
//  b  **  **
//  c
//  d
//  e
//  f
//  code x78
//  0
//  1
//  2
//  3
//  4
//  5 **    **
//  6  **  **
//  7   ****
//  8    **
//  9   ****
//  a  **  **
//  b **    **
//  c
//  d
//  e
//  f
//  code x79
//  0
//  1
//  2
//  3
//  4
//  5 **   **
//  6 **   **
//  7 **   **
//  8 **   **
//  9 **   **
//  a **   **
//  b  ******
//  c      **
//  d     **
//  e *****
//  f
//  code x7a
//  0
//  1
//  2
//  3
//  4
//  5 *******
//  6 **  **
//  7    **
//  8   **
//  9  **
//  a **   **
//  b *******
//  c
//  d
//  e
//  f
//  code x7b
//  0
//  1
//  2     ***
//  3    **
//  4    **
//  5    **
//  6  ***
//  7    **
//  8    **
//  9    **
//  a    **
//  b     ***
//  c
//  d
//  e
//  f
//  code x7c
//  0
//  1
//  2    **
//  3    **
//  4    **
//  5    **
//  6
//  7    **
//  8    **
//  9    **
//  a    **
//  b    **
//  c
//  d
//  e
//  f
//  code x7d
//  0
//  1
//  2  ***
//  3    **
//  4    **
//  5    **
//  6     ***
//  7    **
//  8    **
//  9    **
//  a    **
//  b  ***
//  c
//  d
//  e
//  f
//  code x7e
//  0
//  1
//  2  *** **
//  3 ** ***
//  4
//  5
//  6
//  7
//  8
//  9
//  a
//  b
//  c
//  d
//  e
//  f
//  code x7f
//  0
//  1
//  2
//  3
//  4    *
//  5   ***
//  6  ** **
//  7 **   **
//  8 **   **
//  9 **   **
//  a *******
//  b
//  c
//  d
//  e
//  f
//  addr register to infer block RAM


always @(posedge clk)
   begin : process_1
   addr_reg <= addr;   
   end

assign data = ROM[
TO_INTEGER(addr_reg)]; 

endmodule // module font_rom

